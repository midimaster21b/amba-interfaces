interface asb_if;
   logic agntx;
   logic areqx;
   logic [31:0] ba;
   logic	bclk;
   logic [31:0] bd;
   logic	berror;
   logic	blast;
   logic	blok;
   logic	bnres;
   logic [1:0]	bprot;
   logic [1:0]	bsize;
   logic [1:0]	btran;
   logic	bwait;
   logic	bwrite;
   logic	dselx;

endinterface // asb_if
